(* keep *)
PS7 ps7_stub(
	.DDRARB				('b0),
	.DMA0ACLK			('b0),
	.DMA0DAREADY			('b0),
	.DMA0DRLAST			('b0),
	.DMA0DRTYPE			('b0),
	.DMA0DRVALID			('b0),
	.DMA1ACLK			('b0),
	.DMA1DAREADY			('b0),
	.DMA1DRLAST			('b0),
	.DMA1DRTYPE			('b0),
	.DMA1DRVALID			('b0),
	.DMA2ACLK			('b0),
	.DMA2DAREADY			('b0),
	.DMA2DRLAST			('b0),
	.DMA2DRTYPE			('b0),
	.DMA2DRVALID			('b0),
	.DMA3ACLK			('b0),
	.DMA3DAREADY			('b0),
	.DMA3DRLAST			('b0),
	.DMA3DRTYPE			('b0),
	.DMA3DRVALID			('b0),
	.EMIOCAN0PHYRX			('b0),
	.EMIOCAN1PHYRX			('b0),
	.EMIOENET0EXTINTIN		('b0),
	.EMIOENET0GMIICOL		('b0),
	.EMIOENET0GMIICRS		('b0),
	.EMIOENET0GMIIRXCLK		('b0),
	.EMIOENET0GMIIRXD		('b0),
	.EMIOENET0GMIIRXDV		('b0),
	.EMIOENET0GMIIRXER		('b0),
	.EMIOENET0GMIITXCLK		('b0),
	.EMIOENET0MDIOI			('b0),
	.EMIOENET1EXTINTIN		('b0),
	.EMIOENET1GMIICOL		('b0),
	.EMIOENET1GMIICRS		('b0),
	.EMIOENET1GMIIRXCLK		('b0),
	.EMIOENET1GMIIRXD		('b0),
	.EMIOENET1GMIIRXDV		('b0),
	.EMIOENET1GMIIRXER		('b0),
	.EMIOENET1GMIITXCLK		('b0),
	.EMIOENET1MDIOI			('b0),
	.EMIOGPIOI			('b0),
	.EMIOI2C0SCLI			('b0),
	.EMIOI2C0SDAI			('b0),
	.EMIOI2C1SCLI			('b0),
	.EMIOI2C1SDAI			('b0),
	.EMIOPJTAGTCK			('b0),
	.EMIOPJTAGTDI			('b0),
	.EMIOPJTAGTMS			('b0),
	.EMIOSDIO0CDN			('b0),
	.EMIOSDIO0CLKFB			('b0),
	.EMIOSDIO0CMDI			('b0),
	.EMIOSDIO0DATAI			('b0),
	.EMIOSDIO0WP			('b0),
	.EMIOSDIO1CDN			('b0),
	.EMIOSDIO1CLKFB			('b0),
	.EMIOSDIO1CMDI			('b0),
	.EMIOSDIO1DATAI			('b0),
	.EMIOSDIO1WP			('b0),
	.EMIOSPI0MI			('b0),
	.EMIOSPI0SCLKI			('b0),
	.EMIOSPI0SI			('b0),
	.EMIOSPI0SSIN			('b0),
	.EMIOSPI1MI			('b0),
	.EMIOSPI1SCLKI			('b0),
	.EMIOSPI1SI			('b0),
	.EMIOSPI1SSIN			('b0),
	.EMIOSRAMINTIN			('b0),
	.EMIOTRACECLK			('b0),
	.EMIOTTC0CLKI			('b0),
	.EMIOTTC1CLKI			('b0),
	.EMIOUART0CTSN			('b0),
	.EMIOUART0DCDN			('b0),
	.EMIOUART0DSRN			('b0),
	.EMIOUART0RIN			('b0),
	.EMIOUART0RX			('b0),
	.EMIOUART1CTSN			('b0),
	.EMIOUART1DCDN			('b0),
	.EMIOUART1DSRN			('b0),
	.EMIOUART1RIN			('b0),
	.EMIOUART1RX			('b0),
	.EMIOUSB0VBUSPWRFAULT		('b0),
	.EMIOUSB1VBUSPWRFAULT		('b0),
	.EMIOWDTCLKI			('b0),
	.EVENTEVENTI			('b0),
	.FCLKCLKTRIGN			('b0),
	.FPGAIDLEN			('b0),
	.FTMDTRACEINATID			('b0),
	.FTMDTRACEINCLOCK		('b0),
	.FTMDTRACEINDATA			('b0),
	.FTMDTRACEINVALID		('b0),
	.FTMTF2PDEBUG			('b0),
	.FTMTF2PTRIG			('b0),
	.FTMTP2FTRIGACK			('b0),
	.IRQF2P				('b0),
	.MAXIGP0ACLK			('b0),
	.MAXIGP0ARREADY			('b0),
	.MAXIGP0AWREADY			('b0),
	.MAXIGP0BID			('b0),
	.MAXIGP0BRESP			('b0),
	.MAXIGP0BVALID			('b0),
	.MAXIGP0RDATA			('b0),
	.MAXIGP0RID			('b0),
	.MAXIGP0RLAST			('b0),
	.MAXIGP0RRESP			('b0),
	.MAXIGP0RVALID			('b0),
	.MAXIGP0WREADY			('b0),
	.MAXIGP1ACLK			('b0),
	.MAXIGP1ARREADY			('b0),
	.MAXIGP1AWREADY			('b0),
	.MAXIGP1BID			('b0),
	.MAXIGP1BRESP			('b0),
	.MAXIGP1BVALID			('b0),
	.MAXIGP1RDATA			('b0),
	.MAXIGP1RID			('b0),
	.MAXIGP1RLAST			('b0),
	.MAXIGP1RRESP			('b0),
	.MAXIGP1RVALID			('b0),
	.MAXIGP1WREADY			('b0),
	.SAXIACPACLK			('b0),
	.SAXIACPARADDR			('b0),
	.SAXIACPARBURST			('b0),
	.SAXIACPARCACHE			('b0),
	.SAXIACPARID			('b0),
	.SAXIACPARLEN			('b0),
	.SAXIACPARLOCK			('b0),
	.SAXIACPARPROT			('b0),
	.SAXIACPARQOS			('b0),
	.SAXIACPARSIZE			('b0),
	.SAXIACPARUSER			('b0),
	.SAXIACPARVALID			('b0),
	.SAXIACPAWADDR			('b0),
	.SAXIACPAWBURST			('b0),
	.SAXIACPAWCACHE			('b0),
	.SAXIACPAWID			('b0),
	.SAXIACPAWLEN			('b0),
	.SAXIACPAWLOCK			('b0),
	.SAXIACPAWPROT			('b0),
	.SAXIACPAWQOS			('b0),
	.SAXIACPAWSIZE			('b0),
	.SAXIACPAWUSER			('b0),
	.SAXIACPAWVALID			('b0),
	.SAXIACPBREADY			('b0),
	.SAXIACPRREADY			('b0),
	.SAXIACPWDATA			('b0),
	.SAXIACPWID			('b0),
	.SAXIACPWLAST			('b0),
	.SAXIACPWSTRB			('b0),
	.SAXIACPWVALID			('b0),
	.SAXIGP0ACLK			('b0),
	.SAXIGP0ARADDR			('b0),
	.SAXIGP0ARBURST			('b0),
	.SAXIGP0ARCACHE			('b0),
	.SAXIGP0ARID			('b0),
	.SAXIGP0ARLEN			('b0),
	.SAXIGP0ARLOCK			('b0),
	.SAXIGP0ARPROT			('b0),
	.SAXIGP0ARQOS			('b0),
	.SAXIGP0ARSIZE			('b0),
	.SAXIGP0ARVALID			('b0),
	.SAXIGP0AWADDR			('b0),
	.SAXIGP0AWBURST			('b0),
	.SAXIGP0AWCACHE			('b0),
	.SAXIGP0AWID			('b0),
	.SAXIGP0AWLEN			('b0),
	.SAXIGP0AWLOCK			('b0),
	.SAXIGP0AWPROT			('b0),
	.SAXIGP0AWQOS			('b0),
	.SAXIGP0AWSIZE			('b0),
	.SAXIGP0AWVALID			('b0),
	.SAXIGP0BREADY			('b0),
	.SAXIGP0RREADY			('b0),
	.SAXIGP0WDATA			('b0),
	.SAXIGP0WID			('b0),
	.SAXIGP0WLAST			('b0),
	.SAXIGP0WSTRB			('b0),
	.SAXIGP0WVALID			('b0),
	.SAXIGP1ACLK			('b0),
	.SAXIGP1ARADDR			('b0),
	.SAXIGP1ARBURST			('b0),
	.SAXIGP1ARCACHE			('b0),
	.SAXIGP1ARID			('b0),
	.SAXIGP1ARLEN			('b0),
	.SAXIGP1ARLOCK			('b0),
	.SAXIGP1ARPROT			('b0),
	.SAXIGP1ARQOS			('b0),
	.SAXIGP1ARSIZE			('b0),
	.SAXIGP1ARVALID			('b0),
	.SAXIGP1AWADDR			('b0),
	.SAXIGP1AWBURST			('b0),
	.SAXIGP1AWCACHE			('b0),
	.SAXIGP1AWID			('b0),
	.SAXIGP1AWLEN			('b0),
	.SAXIGP1AWLOCK			('b0),
	.SAXIGP1AWPROT			('b0),
	.SAXIGP1AWQOS			('b0),
	.SAXIGP1AWSIZE			('b0),
	.SAXIGP1AWVALID			('b0),
	.SAXIGP1BREADY			('b0),
	.SAXIGP1RREADY			('b0),
	.SAXIGP1WDATA			('b0),
	.SAXIGP1WID			('b0),
	.SAXIGP1WLAST			('b0),
	.SAXIGP1WSTRB			('b0),
	.SAXIGP1WVALID			('b0),
	.SAXIHP0ACLK			('b0),
	.SAXIHP0ARADDR			('b0),
	.SAXIHP0ARBURST			('b0),
	.SAXIHP0ARCACHE			('b0),
	.SAXIHP0ARID			('b0),
	.SAXIHP0ARLEN			('b0),
	.SAXIHP0ARLOCK			('b0),
	.SAXIHP0ARPROT			('b0),
	.SAXIHP0ARQOS			('b0),
	.SAXIHP0ARSIZE			('b0),
	.SAXIHP0ARVALID			('b0),
	.SAXIHP0AWADDR			('b0),
	.SAXIHP0AWBURST			('b0),
	.SAXIHP0AWCACHE			('b0),
	.SAXIHP0AWID			('b0),
	.SAXIHP0AWLEN			('b0),
	.SAXIHP0AWLOCK			('b0),
	.SAXIHP0AWPROT			('b0),
	.SAXIHP0AWQOS			('b0),
	.SAXIHP0AWSIZE			('b0),
	.SAXIHP0AWVALID			('b0),
	.SAXIHP0BREADY			('b0),
	.SAXIHP0RDISSUECAP1EN		('b0),
	.SAXIHP0RREADY			('b0),
	.SAXIHP0WDATA			('b0),
	.SAXIHP0WID			('b0),
	.SAXIHP0WLAST			('b0),
	.SAXIHP0WRISSUECAP1EN		('b0),
	.SAXIHP0WSTRB			('b0),
	.SAXIHP0WVALID			('b0),
	.SAXIHP1ACLK			('b0),
	.SAXIHP1ARADDR			('b0),
	.SAXIHP1ARBURST			('b0),
	.SAXIHP1ARCACHE			('b0),
	.SAXIHP1ARID			('b0),
	.SAXIHP1ARLEN			('b0),
	.SAXIHP1ARLOCK			('b0),
	.SAXIHP1ARPROT			('b0),
	.SAXIHP1ARQOS			('b0),
	.SAXIHP1ARSIZE			('b0),
	.SAXIHP1ARVALID			('b0),
	.SAXIHP1AWADDR			('b0),
	.SAXIHP1AWBURST			('b0),
	.SAXIHP1AWCACHE			('b0),
	.SAXIHP1AWID			('b0),
	.SAXIHP1AWLEN			('b0),
	.SAXIHP1AWLOCK			('b0),
	.SAXIHP1AWPROT			('b0),
	.SAXIHP1AWQOS			('b0),
	.SAXIHP1AWSIZE			('b0),
	.SAXIHP1AWVALID			('b0),
	.SAXIHP1BREADY			('b0),
	.SAXIHP1RDISSUECAP1EN		('b0),
	.SAXIHP1RREADY			('b0),
	.SAXIHP1WDATA			('b0),
	.SAXIHP1WID			('b0),
	.SAXIHP1WLAST			('b0),
	.SAXIHP1WRISSUECAP1EN		('b0),
	.SAXIHP1WSTRB			('b0),
	.SAXIHP1WVALID			('b0),
	.SAXIHP2ACLK			('b0),
	.SAXIHP2ARADDR			('b0),
	.SAXIHP2ARBURST			('b0),
	.SAXIHP2ARCACHE			('b0),
	.SAXIHP2ARID			('b0),
	.SAXIHP2ARLEN			('b0),
	.SAXIHP2ARLOCK			('b0),
	.SAXIHP2ARPROT			('b0),
	.SAXIHP2ARQOS			('b0),
	.SAXIHP2ARSIZE			('b0),
	.SAXIHP2ARVALID			('b0),
	.SAXIHP2AWADDR			('b0),
	.SAXIHP2AWBURST			('b0),
	.SAXIHP2AWCACHE			('b0),
	.SAXIHP2AWID			('b0),
	.SAXIHP2AWLEN			('b0),
	.SAXIHP2AWLOCK			('b0),
	.SAXIHP2AWPROT			('b0),
	.SAXIHP2AWQOS			('b0),
	.SAXIHP2AWSIZE			('b0),
	.SAXIHP2AWVALID			('b0),
	.SAXIHP2BREADY			('b0),
	.SAXIHP2RDISSUECAP1EN		('b0),
	.SAXIHP2RREADY			('b0),
	.SAXIHP2WDATA			('b0),
	.SAXIHP2WID			('b0),
	.SAXIHP2WLAST			('b0),
	.SAXIHP2WRISSUECAP1EN		('b0),
	.SAXIHP2WSTRB			('b0),
	.SAXIHP2WVALID			('b0),
	.SAXIHP3ACLK			('b0),
	.SAXIHP3ARADDR			('b0),
	.SAXIHP3ARBURST			('b0),
	.SAXIHP3ARCACHE			('b0),
	.SAXIHP3ARID			('b0),
	.SAXIHP3ARLEN			('b0),
	.SAXIHP3ARLOCK			('b0),
	.SAXIHP3ARPROT			('b0),
	.SAXIHP3ARQOS			('b0),
	.SAXIHP3ARSIZE			('b0),
	.SAXIHP3ARVALID			('b0),
	.SAXIHP3AWADDR			('b0),
	.SAXIHP3AWBURST			('b0),
	.SAXIHP3AWCACHE			('b0),
	.SAXIHP3AWID			('b0),
	.SAXIHP3AWLEN			('b0),
	.SAXIHP3AWLOCK			('b0),
	.SAXIHP3AWPROT			('b0),
	.SAXIHP3AWQOS			('b0),
	.SAXIHP3AWSIZE			('b0),
	.SAXIHP3AWVALID			('b0),
	.SAXIHP3BREADY			('b0),
	.SAXIHP3RDISSUECAP1EN		('b0),
	.SAXIHP3RREADY			('b0),
	.SAXIHP3WDATA			('b0),
	.SAXIHP3WID			('b0),
	.SAXIHP3WLAST			('b0),
	.SAXIHP3WRISSUECAP1EN		('b0),
	.SAXIHP3WSTRB			('b0),
	.SAXIHP3WVALID			('b0)
);
