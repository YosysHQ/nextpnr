module top(output o, output o2);

assign o = 1'b0;
assign o2 = 1'b1;

endmodule
