module top(input i0, input i1, output o);

assign o = i0 | i1;

endmodule
