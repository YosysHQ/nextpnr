module top(output o, output o2, output o3, output o4);

assign o = 1'b0;
assign o2 = 1'b1;
assign o3 = 1'b0;
assign o4 = 1'b1;

endmodule
